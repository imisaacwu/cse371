/* Arbitrary ASM chart implementation to examine output timings */
module hw3p3 (clk, reset, X, Ya, Yb, Yc, Z1, Z2);
	
	// for you to implement
	
endmodule  // hw3p3
