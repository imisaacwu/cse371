/* Testbench for Homework 3 Problem 3 */
module hw3p3_tb ();
	
	// for you to implement
	
	hw3p3 dut (.*);
	
	initial begin
		
		// for you to implement
		
	end  // initial
	
endmodule  // hw3p3_tb
